`include"MCS_dv05_subtractor_dut.sv"
`include"MCS_dv05_subtractor_transaction1.sv"
`include"MCS_dv05_subtractor_generator2.sv"
`include"MCS_dv05_subtractor_interface.sv"
`include"MCS_dv05_subtractor_driver3.sv"
`include"MCS_dv05_subtractor_input_monitor_checker.sv"
`include"MCS_dv05_subtractor_op_monitor_from_dut.sv"
`include"MCS_dv05_subtractor_scoreboard_comparator.sv"
`include"MCS_dv05_subtractor_environment.sv"
`include"test.sv"
`include"MCS_dv05_subtractor_top.sv"
