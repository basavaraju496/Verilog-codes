`include"1_transaction.sv"

`include"2_generator.sv"   // do var

`include"3_interface.sv"   // do var with delays

`include"4_driver.sv"   // do var with blocking and non blocking

`include"5_checker.sv"   // do var with blocking and non blocking

`include"6_dut_monitor.sv"   // do var with blocking and non blocking

`include"7_score_board.sv"   // do var with blocking and non blocking








