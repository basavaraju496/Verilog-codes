class driver;



mailbox hmb1;

transaction ht2;

function new(,mailbox mb1)
		hmb1=mb1;
		endfunction







endclass
